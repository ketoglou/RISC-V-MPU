-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.0 Build 156 04/24/2013 SJ Web Edition"
-- CREATED		"Sun Feb 07 20:49:44 2021"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY RISCV_CPU IS 
	PORT
	(
		CLK :  IN  STD_LOGIC;
		CLEAR :  IN  STD_LOGIC;
		PIN1_IN :  IN  STD_LOGIC;
		MEM_WR :  IN  STD_LOGIC;
		DATAWR :  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		PIN2_OUT :  OUT  STD_LOGIC;
		PIN3_OUT :  OUT  STD_LOGIC;
		PIN4_OUT :  OUT  STD_LOGIC;
		PIN5_OUT :  OUT  STD_LOGIC
	);
END RISCV_CPU;

ARCHITECTURE bdf_type OF RISCV_CPU IS 

COMPONENT instruction_memory
	PORT(MEM_WR : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 ADDRESS_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA_WR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT mux2_32
	PORT(SEL : IN STD_LOGIC;
		 D0 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 D1 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Y : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT cla_32_pc_add
	PORT(A : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 B : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 S : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT register_rd_csr
	PORT(CLK : IN STD_LOGIC;
		 CLR : IN STD_LOGIC;
		 CSR : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
		 RD : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 CSR_O : OUT STD_LOGIC_VECTOR(11 DOWNTO 0);
		 RD_O : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
	);
END COMPONENT;

COMPONENT register_32
	PORT(CLK : IN STD_LOGIC;
		 CLR : IN STD_LOGIC;
		 HOLD : IN STD_LOGIC;
		 D_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 D_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT jump_branch_exception
	PORT(NEW_PC : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 JB_EXCEPTION : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT exp_int_handler
	PORT(MRET_EN : IN STD_LOGIC;
		 OP_EXP : IN STD_LOGIC;
		 JB_EXP : IN STD_LOGIC;
		 INT_EXTERNAL : IN STD_LOGIC;
		 CSR_WR : IN STD_LOGIC;
		 EXP_INT_EN_RETURN : IN STD_LOGIC;
		 CLR : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 CSR_ADDRESS : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
		 CSR_ADDRESS_WR : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
		 CSR_DATA_WR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 INVALID_ADDRESS : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 INVALID_INST : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
		 PC : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 EXP_INT_EN : OUT STD_LOGIC;
		 CSR_DATA : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 EXP_INT_PC : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT mux8_1
	PORT(D0 : IN STD_LOGIC;
		 D1 : IN STD_LOGIC;
		 D2 : IN STD_LOGIC;
		 D3 : IN STD_LOGIC;
		 D4 : IN STD_LOGIC;
		 D5 : IN STD_LOGIC;
		 D6 : IN STD_LOGIC;
		 D7 : IN STD_LOGIC;
		 SEL : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 Y : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT data_hazard_unit
	PORT(OPCODE : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		 RD_ID_EX : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 RS1_IF_ID : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 RS2_IF_ID : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 WR_ID_EX : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 DH_EN : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT registers_id
	PORT(CLR : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 CSR : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
		 RD : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 RS1 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 RS2 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 CSR_O : OUT STD_LOGIC_VECTOR(11 DOWNTO 0);
		 RD_O : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
		 RS1_O : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
		 RS2_O : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
	);
END COMPONENT;

COMPONENT data_memory
	PORT(MEM_WR : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 ADDRESS_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA_WR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 MEM_OP : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 DATA_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 EXP_PINS : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT x_registers
	PORT(WR : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 DATA_WRITE : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 RD : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 RS1 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 RS2 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 DATA1 : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA2 : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT forwarding_unit
	PORT(WB_EX_MEM : IN STD_LOGIC;
		 WB_MEM_WB : IN STD_LOGIC;
		 EN_IMM : IN STD_LOGIC;
		 RD_EX_MEM : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 RD_MEM_WB : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 RS1_ID : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 RS1_ID_EX : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 RS2_ID : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 RS2_ID_EX : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 FORWARD_ID1 : OUT STD_LOGIC;
		 FORWARD_ID2 : OUT STD_LOGIC;
		 FORWARD_1 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		 FORWARD_2 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	);
END COMPONENT;

COMPONENT mux4_32
	PORT(D0 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 D1 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 D2 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 D3 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 SEL : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 Y : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT register_array_3
	PORT(CLR : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 HOLD : IN STD_LOGIC;
		 DATA1_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA2_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA3_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA1_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA2_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA3_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT register_array_6
	PORT(CLR : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 DATA1_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA2_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA3_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA4_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA5_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA6_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA1_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA2_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA3_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA4_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA5_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA6_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT not_unit
	PORT(NOT_ENABLE : IN STD_LOGIC;
		 DATA_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT register_array_7
	PORT(CLR : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 DATA1_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA2_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA3_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA4_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA5_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA6_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA7_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA1_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA2_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA3_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA4_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA5_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA6_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA7_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT sign_extension
	PORT(INST : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 IMMEDIATE : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT mux8_32
	PORT(D0 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 D1 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 D2 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 D3 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 D4 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 D5 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 D6 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 D7 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 SEL : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 Y : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT control_unit
	PORT(FUNCT3 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 FUNCT7 : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		 OPCODE : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		 CSR_WB : OUT STD_LOGIC;
		 WB : OUT STD_LOGIC;
		 BRANCH : OUT STD_LOGIC;
		 MEM_WR : OUT STD_LOGIC;
		 EX1 : OUT STD_LOGIC;
		 EN_IMM : OUT STD_LOGIC;
		 C1 : OUT STD_LOGIC;
		 C2 : OUT STD_LOGIC;
		 NE1 : OUT STD_LOGIC;
		 NE2 : OUT STD_LOGIC;
		 OP_EXP : OUT STD_LOGIC;
		 MRET_EN : OUT STD_LOGIC;
		 ALU_OP : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 WR : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
	);
END COMPONENT;

COMPONENT pip_reg_id_exe
	PORT(CSR_WB : IN STD_LOGIC;
		 WB : IN STD_LOGIC;
		 BRANCH : IN STD_LOGIC;
		 MEM_WR : IN STD_LOGIC;
		 EX1 : IN STD_LOGIC;
		 EN_IMM : IN STD_LOGIC;
		 C1 : IN STD_LOGIC;
		 C2 : IN STD_LOGIC;
		 NE1 : IN STD_LOGIC;
		 NE2 : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 CLR : IN STD_LOGIC;
		 ALU_OP : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 FUNCT3 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 WR : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 CSR_WB_O : OUT STD_LOGIC;
		 WB_O : OUT STD_LOGIC;
		 BRANCH_O : OUT STD_LOGIC;
		 MEM_WR_O : OUT STD_LOGIC;
		 EX1_O : OUT STD_LOGIC;
		 EN_IMM_O : OUT STD_LOGIC;
		 C1_O : OUT STD_LOGIC;
		 C2_O : OUT STD_LOGIC;
		 NE1_O : OUT STD_LOGIC;
		 NE2_O : OUT STD_LOGIC;
		 ALU_OP_O : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 FUNCT3_O : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		 WR_O : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
	);
END COMPONENT;

COMPONENT pip_reg_exe_mem
	PORT(CSR_WB : IN STD_LOGIC;
		 WB : IN STD_LOGIC;
		 BRANCH : IN STD_LOGIC;
		 MEM_WR : IN STD_LOGIC;
		 ZERO : IN STD_LOGIC;
		 LESS_THAN_SIGNED : IN STD_LOGIC;
		 LESS_THAN_UNSIGNED : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 CLR : IN STD_LOGIC;
		 FUNCT3 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 WR : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 CSR_WB_O : OUT STD_LOGIC;
		 WB_O : OUT STD_LOGIC;
		 BRANCH_O : OUT STD_LOGIC;
		 ZERO_O : OUT STD_LOGIC;
		 LESS_THAN_SIGNED_O : OUT STD_LOGIC;
		 LESS_THAN_UNSIGNED_O : OUT STD_LOGIC;
		 MEM_WR_O : OUT STD_LOGIC;
		 FUNCT3_O : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		 WR_O : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
	);
END COMPONENT;

COMPONENT pip_reg_mem_wb
	PORT(CSR_WB : IN STD_LOGIC;
		 WB : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 CLR : IN STD_LOGIC;
		 WR : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 CSR_WB_O : OUT STD_LOGIC;
		 WB_O : OUT STD_LOGIC;
		 WR_O : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
	);
END COMPONENT;

COMPONENT flag_reg
	PORT(FLAG_IN : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 CLR : IN STD_LOGIC;
		 FLAG_OUT : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT cla_32_add_1
	PORT(A : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 S : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT alu
	PORT(DATAIN_1 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATAIN_2 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 OP : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 ZERO : OUT STD_LOGIC;
		 LESS_THAN_SIGNED : OUT STD_LOGIC;
		 LESS_THAN_UNSIGNED : OUT STD_LOGIC;
		 DATA_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	ALU_OP :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	C1_O :  STD_LOGIC;
SIGNAL	C2_O :  STD_LOGIC;
SIGNAL	CSR_DATA :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	CSR_WB_O :  STD_LOGIC;
SIGNAL	DATA1 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	DATA2 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	DH_EN :  STD_LOGIC;
SIGNAL	EN_IMM_O :  STD_LOGIC;
SIGNAL	EX1_O :  STD_LOGIC;
SIGNAL	EXP_INT_EN :  STD_LOGIC;
SIGNAL	EXP_INT_PC :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	EXP_INT_RETURN :  STD_LOGIC;
SIGNAL	EXP_PINS :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	FLUSH :  STD_LOGIC;
SIGNAL	FLUSH_BJ :  STD_LOGIC;
SIGNAL	FORWARD_1 :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	FORWARD_2 :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	FORWARD_ID1 :  STD_LOGIC;
SIGNAL	FORWARD_ID2 :  STD_LOGIC;
SIGNAL	FUNCT3 :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	ID :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	IMM :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	INT_EXTERNAL :  STD_LOGIC;
SIGNAL	INV_ADDRESS :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	JB_EXP :  STD_LOGIC;
SIGNAL	MEM_WR_O :  STD_LOGIC;
SIGNAL	MRET_EN :  STD_LOGIC;
SIGNAL	NE1_O :  STD_LOGIC;
SIGNAL	NE2_O :  STD_LOGIC;
SIGNAL	OP_EXP :  STD_LOGIC;
SIGNAL	PC :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	PC_4 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	PC_ID :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	RD_O :  STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL	WB_O :  STD_LOGIC;
SIGNAL	WR2_IE :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	WR_O :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_100 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_101 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC_VECTOR(11 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC_VECTOR(11 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_102 :  STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_103 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_104 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC_VECTOR(11 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_105 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_106 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_107 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_108 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_109 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_110 :  STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_111 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_55 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_58 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_59 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_60 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_61 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_62 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_64 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_65 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_66 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_67 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_68 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_69 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_70 :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_71 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_72 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_73 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_74 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_75 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_76 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_77 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_78 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_79 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_80 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_81 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_82 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_83 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_84 :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_87 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_88 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_89 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_90 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_91 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_92 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_93 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_94 :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_95 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_96 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_98 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_99 :  STD_LOGIC_VECTOR(31 DOWNTO 0);


BEGIN 



b2v_inst : instruction_memory
PORT MAP(MEM_WR => MEM_WR,
		 CLK => CLK,
		 ADDRESS_IN => SYNTHESIZED_WIRE_100,
		 DATA_WR => DATAWR,
		 DATA_OUT => SYNTHESIZED_WIRE_41);


b2v_inst1 : mux2_32
PORT MAP(SEL => FLUSH_BJ,
		 D0 => SYNTHESIZED_WIRE_101,
		 D1 => INV_ADDRESS,
		 Y => SYNTHESIZED_WIRE_33);


b2v_inst10 : cla_32_pc_add
PORT MAP(A => IMM,
		 B => SYNTHESIZED_WIRE_2,
		 S => SYNTHESIZED_WIRE_56);


b2v_inst11 : register_rd_csr
PORT MAP(CLK => CLK,
		 CLR => CLEAR,
		 CSR => SYNTHESIZED_WIRE_3,
		 RD => RD_O,
		 CSR_O => SYNTHESIZED_WIRE_4,
		 RD_O => SYNTHESIZED_WIRE_102);


b2v_inst12 : register_rd_csr
PORT MAP(CLK => CLK,
		 CLR => CLEAR,
		 CSR => SYNTHESIZED_WIRE_4,
		 RD => SYNTHESIZED_WIRE_102,
		 CSR_O => SYNTHESIZED_WIRE_12,
		 RD_O => SYNTHESIZED_WIRE_110);


b2v_inst13 : register_32
PORT MAP(CLK => CLK,
		 CLR => CLEAR,
		 HOLD => SYNTHESIZED_WIRE_6,
		 D_IN => SYNTHESIZED_WIRE_7,
		 D_OUT => SYNTHESIZED_WIRE_100);


b2v_inst14 : mux2_32
PORT MAP(SEL => FORWARD_ID1,
		 D0 => SYNTHESIZED_WIRE_8,
		 D1 => SYNTHESIZED_WIRE_103,
		 Y => SYNTHESIZED_WIRE_43);


b2v_inst15 : jump_branch_exception
PORT MAP(NEW_PC => INV_ADDRESS,
		 JB_EXCEPTION => SYNTHESIZED_WIRE_10);


JB_EXP <= FLUSH_BJ AND SYNTHESIZED_WIRE_10;


b2v_inst17 : exp_int_handler
PORT MAP(MRET_EN => MRET_EN,
		 OP_EXP => OP_EXP,
		 JB_EXP => JB_EXP,
		 INT_EXTERNAL => INT_EXTERNAL,
		 CSR_WR => SYNTHESIZED_WIRE_104,
		 EXP_INT_EN_RETURN => EXP_INT_RETURN,
		 CLR => CLEAR,
		 CLK => CLK,
		 CSR_ADDRESS => ID(31 DOWNTO 20),
		 CSR_ADDRESS_WR => SYNTHESIZED_WIRE_12,
		 CSR_DATA_WR => SYNTHESIZED_WIRE_105,
		 INVALID_ADDRESS => INV_ADDRESS,
		 INVALID_INST => ID(19 DOWNTO 0),
		 PC => PC_ID,
		 EXP_INT_EN => EXP_INT_EN,
		 CSR_DATA => SYNTHESIZED_WIRE_46,
		 EXP_INT_PC => EXP_INT_PC);


b2v_inst18 : mux8_1
PORT MAP(D0 => SYNTHESIZED_WIRE_106,
		 D1 => SYNTHESIZED_WIRE_15,
		 D2 => '0',
		 D3 => '0',
		 D4 => SYNTHESIZED_WIRE_107,
		 D5 => SYNTHESIZED_WIRE_17,
		 D6 => SYNTHESIZED_WIRE_108,
		 D7 => SYNTHESIZED_WIRE_19,
		 SEL => FUNCT3,
		 Y => SYNTHESIZED_WIRE_72);


b2v_inst19 : data_hazard_unit
PORT MAP(OPCODE => ID(6 DOWNTO 0),
		 RD_ID_EX => RD_O,
		 RS1_IF_ID => ID(19 DOWNTO 15),
		 RS2_IF_ID => ID(24 DOWNTO 20),
		 WR_ID_EX => WR2_IE,
		 DH_EN => DH_EN);


b2v_inst2 : registers_id
PORT MAP(CLR => FLUSH,
		 CLK => CLK,
		 CSR => ID(31 DOWNTO 20),
		 RD => ID(11 DOWNTO 7),
		 RS1 => ID(19 DOWNTO 15),
		 RS2 => ID(24 DOWNTO 20),
		 CSR_O => SYNTHESIZED_WIRE_3,
		 RD_O => RD_O,
		 RS1_O => SYNTHESIZED_WIRE_30,
		 RS2_O => SYNTHESIZED_WIRE_31);


SYNTHESIZED_WIRE_15 <= NOT(SYNTHESIZED_WIRE_106);



SYNTHESIZED_WIRE_38 <= FLUSH_BJ OR MRET_EN OR CLEAR;


b2v_inst22 : data_memory
PORT MAP(MEM_WR => MEM_WR_O,
		 CLK => CLK,
		 ADDRESS_IN => INV_ADDRESS,
		 DATA_WR => SYNTHESIZED_WIRE_21,
		 MEM_OP => FUNCT3,
		 DATA_OUT => SYNTHESIZED_WIRE_62,
		 EXP_PINS => EXP_PINS);


b2v_inst24 : mux2_32
PORT MAP(SEL => FORWARD_ID2,
		 D0 => SYNTHESIZED_WIRE_22,
		 D1 => SYNTHESIZED_WIRE_103,
		 Y => SYNTHESIZED_WIRE_44);


b2v_inst25 : x_registers
PORT MAP(WR => SYNTHESIZED_WIRE_109,
		 CLK => CLK,
		 DATA_WRITE => SYNTHESIZED_WIRE_103,
		 RD => SYNTHESIZED_WIRE_110,
		 RS1 => ID(19 DOWNTO 15),
		 RS2 => ID(24 DOWNTO 20),
		 DATA1 => SYNTHESIZED_WIRE_8,
		 DATA2 => SYNTHESIZED_WIRE_22);


b2v_inst26 : forwarding_unit
PORT MAP(WB_EX_MEM => WB_O,
		 WB_MEM_WB => SYNTHESIZED_WIRE_109,
		 EN_IMM => EN_IMM_O,
		 RD_EX_MEM => SYNTHESIZED_WIRE_102,
		 RD_MEM_WB => SYNTHESIZED_WIRE_110,
		 RS1_ID => ID(19 DOWNTO 15),
		 RS1_ID_EX => SYNTHESIZED_WIRE_30,
		 RS2_ID => ID(24 DOWNTO 20),
		 RS2_ID_EX => SYNTHESIZED_WIRE_31,
		 FORWARD_ID1 => FORWARD_ID1,
		 FORWARD_ID2 => FORWARD_ID2,
		 FORWARD_1 => FORWARD_1,
		 FORWARD_2 => FORWARD_2);


FLUSH <= CLEAR OR FLUSH_BJ OR DH_EN;


SYNTHESIZED_WIRE_6 <= SYNTHESIZED_WIRE_32 AND DH_EN;


b2v_inst3 : mux2_32
PORT MAP(SEL => EXP_INT_EN,
		 D0 => SYNTHESIZED_WIRE_33,
		 D1 => EXP_INT_PC,
		 Y => SYNTHESIZED_WIRE_7);


SYNTHESIZED_WIRE_32 <= NOT(FLUSH_BJ);



b2v_inst33 : mux4_32
PORT MAP(D0 => DATA2,
		 D1 => SYNTHESIZED_WIRE_111,
		 D2 => SYNTHESIZED_WIRE_105,
		 D3 => IMM,
		 SEL => FORWARD_2,
		 Y => SYNTHESIZED_WIRE_55);


b2v_inst34 : mux4_32
PORT MAP(D0 => DATA1,
		 D1 => SYNTHESIZED_WIRE_111,
		 D2 => SYNTHESIZED_WIRE_105,
		 D3 => x"00000000",
		 SEL => FORWARD_1,
		 Y => SYNTHESIZED_WIRE_51);


b2v_inst35 : register_array_3
PORT MAP(CLR => SYNTHESIZED_WIRE_38,
		 CLK => CLK,
		 HOLD => DH_EN,
		 DATA1_IN => SYNTHESIZED_WIRE_101,
		 DATA2_IN => SYNTHESIZED_WIRE_100,
		 DATA3_IN => SYNTHESIZED_WIRE_41,
		 DATA1_OUT => SYNTHESIZED_WIRE_42,
		 DATA2_OUT => PC_ID,
		 DATA3_OUT => ID);


b2v_inst36 : register_array_6
PORT MAP(CLR => FLUSH,
		 CLK => CLK,
		 DATA1_IN => SYNTHESIZED_WIRE_42,
		 DATA2_IN => PC_ID,
		 DATA3_IN => SYNTHESIZED_WIRE_43,
		 DATA4_IN => SYNTHESIZED_WIRE_44,
		 DATA5_IN => SYNTHESIZED_WIRE_45,
		 DATA6_IN => SYNTHESIZED_WIRE_46,
		 DATA1_OUT => PC_4,
		 DATA2_OUT => PC,
		 DATA3_OUT => DATA1,
		 DATA4_OUT => DATA2,
		 DATA5_OUT => IMM,
		 DATA6_OUT => CSR_DATA);


b2v_inst38 : mux2_32
PORT MAP(SEL => SYNTHESIZED_WIRE_104,
		 D0 => SYNTHESIZED_WIRE_105,
		 D1 => SYNTHESIZED_WIRE_49,
		 Y => SYNTHESIZED_WIRE_103);


b2v_inst4 : mux2_32
PORT MAP(SEL => EX1_O,
		 D0 => PC,
		 D1 => DATA1,
		 Y => SYNTHESIZED_WIRE_2);


b2v_inst43 : mux2_32
PORT MAP(SEL => C1_O,
		 D0 => SYNTHESIZED_WIRE_50,
		 D1 => CSR_DATA,
		 Y => SYNTHESIZED_WIRE_98);


b2v_inst44 : not_unit
PORT MAP(NOT_ENABLE => NE1_O,
		 DATA_IN => SYNTHESIZED_WIRE_51,
		 DATA_OUT => SYNTHESIZED_WIRE_50);


b2v_inst45 : mux2_32
PORT MAP(SEL => C2_O,
		 D0 => SYNTHESIZED_WIRE_52,
		 D1 => CSR_DATA,
		 Y => SYNTHESIZED_WIRE_99);


FLUSH_BJ <= SYNTHESIZED_WIRE_53 OR SYNTHESIZED_WIRE_54;


b2v_inst48 : not_unit
PORT MAP(NOT_ENABLE => NE2_O,
		 DATA_IN => SYNTHESIZED_WIRE_55,
		 DATA_OUT => SYNTHESIZED_WIRE_52);


b2v_inst49 : register_array_7
PORT MAP(CLR => CLEAR,
		 CLK => CLK,
		 DATA1_IN => SYNTHESIZED_WIRE_56,
		 DATA2_IN => PC_4,
		 DATA3_IN => IMM,
		 DATA4_IN => DATA1,
		 DATA5_IN => CSR_DATA,
		 DATA6_IN => DATA2,
		 DATA7_IN => SYNTHESIZED_WIRE_57,
		 DATA1_OUT => INV_ADDRESS,
		 DATA2_OUT => SYNTHESIZED_WIRE_58,
		 DATA3_OUT => SYNTHESIZED_WIRE_59,
		 DATA4_OUT => SYNTHESIZED_WIRE_60,
		 DATA5_OUT => SYNTHESIZED_WIRE_61,
		 DATA6_OUT => SYNTHESIZED_WIRE_21,
		 DATA7_OUT => SYNTHESIZED_WIRE_111);


b2v_inst5 : sign_extension
PORT MAP(INST => ID,
		 IMMEDIATE => SYNTHESIZED_WIRE_45);


b2v_inst51 : register_array_7
PORT MAP(CLR => CLEAR,
		 CLK => CLK,
		 DATA1_IN => INV_ADDRESS,
		 DATA2_IN => SYNTHESIZED_WIRE_58,
		 DATA3_IN => SYNTHESIZED_WIRE_59,
		 DATA4_IN => SYNTHESIZED_WIRE_60,
		 DATA5_IN => SYNTHESIZED_WIRE_61,
		 DATA6_IN => SYNTHESIZED_WIRE_62,
		 DATA7_IN => SYNTHESIZED_WIRE_111,
		 DATA1_OUT => SYNTHESIZED_WIRE_64,
		 DATA2_OUT => SYNTHESIZED_WIRE_65,
		 DATA3_OUT => SYNTHESIZED_WIRE_66,
		 DATA4_OUT => SYNTHESIZED_WIRE_67,
		 DATA5_OUT => SYNTHESIZED_WIRE_49,
		 DATA6_OUT => SYNTHESIZED_WIRE_68,
		 DATA7_OUT => SYNTHESIZED_WIRE_69);


b2v_inst52 : mux8_32
PORT MAP(D0 => SYNTHESIZED_WIRE_64,
		 D1 => SYNTHESIZED_WIRE_65,
		 D2 => SYNTHESIZED_WIRE_66,
		 D3 => SYNTHESIZED_WIRE_67,
		 D4 => SYNTHESIZED_WIRE_68,
		 D5 => SYNTHESIZED_WIRE_69,
		 D6 => x"00000000",
		 D7 => x"00000000",
		 SEL => SYNTHESIZED_WIRE_70,
		 Y => SYNTHESIZED_WIRE_105);


b2v_inst53 : control_unit
PORT MAP(FUNCT3 => ID(14 DOWNTO 12),
		 FUNCT7 => ID(31 DOWNTO 25),
		 OPCODE => ID(6 DOWNTO 0),
		 CSR_WB => SYNTHESIZED_WIRE_73,
		 WB => SYNTHESIZED_WIRE_74,
		 BRANCH => SYNTHESIZED_WIRE_75,
		 MEM_WR => SYNTHESIZED_WIRE_76,
		 EX1 => SYNTHESIZED_WIRE_77,
		 EN_IMM => SYNTHESIZED_WIRE_78,
		 C1 => SYNTHESIZED_WIRE_79,
		 C2 => SYNTHESIZED_WIRE_80,
		 NE1 => SYNTHESIZED_WIRE_81,
		 NE2 => SYNTHESIZED_WIRE_82,
		 OP_EXP => OP_EXP,
		 MRET_EN => MRET_EN,
		 ALU_OP => SYNTHESIZED_WIRE_83,
		 WR => SYNTHESIZED_WIRE_84);


SYNTHESIZED_WIRE_54 <= SYNTHESIZED_WIRE_71 AND SYNTHESIZED_WIRE_72;


b2v_inst55 : pip_reg_id_exe
PORT MAP(CSR_WB => SYNTHESIZED_WIRE_73,
		 WB => SYNTHESIZED_WIRE_74,
		 BRANCH => SYNTHESIZED_WIRE_75,
		 MEM_WR => SYNTHESIZED_WIRE_76,
		 EX1 => SYNTHESIZED_WIRE_77,
		 EN_IMM => SYNTHESIZED_WIRE_78,
		 C1 => SYNTHESIZED_WIRE_79,
		 C2 => SYNTHESIZED_WIRE_80,
		 NE1 => SYNTHESIZED_WIRE_81,
		 NE2 => SYNTHESIZED_WIRE_82,
		 CLK => CLK,
		 CLR => FLUSH,
		 ALU_OP => SYNTHESIZED_WIRE_83,
		 FUNCT3 => ID(14 DOWNTO 12),
		 WR => SYNTHESIZED_WIRE_84,
		 CSR_WB_O => SYNTHESIZED_WIRE_87,
		 WB_O => SYNTHESIZED_WIRE_88,
		 BRANCH_O => SYNTHESIZED_WIRE_89,
		 MEM_WR_O => SYNTHESIZED_WIRE_90,
		 EX1_O => EX1_O,
		 EN_IMM_O => EN_IMM_O,
		 C1_O => C1_O,
		 C2_O => C2_O,
		 NE1_O => NE1_O,
		 NE2_O => NE2_O,
		 ALU_OP_O => ALU_OP,
		 FUNCT3_O => SYNTHESIZED_WIRE_94,
		 WR_O => WR2_IE);


SYNTHESIZED_WIRE_17 <= NOT(SYNTHESIZED_WIRE_107);



SYNTHESIZED_WIRE_19 <= NOT(SYNTHESIZED_WIRE_108);



b2v_inst58 : pip_reg_exe_mem
PORT MAP(CSR_WB => SYNTHESIZED_WIRE_87,
		 WB => SYNTHESIZED_WIRE_88,
		 BRANCH => SYNTHESIZED_WIRE_89,
		 MEM_WR => SYNTHESIZED_WIRE_90,
		 ZERO => SYNTHESIZED_WIRE_91,
		 LESS_THAN_SIGNED => SYNTHESIZED_WIRE_92,
		 LESS_THAN_UNSIGNED => SYNTHESIZED_WIRE_93,
		 CLK => CLK,
		 CLR => CLEAR,
		 FUNCT3 => SYNTHESIZED_WIRE_94,
		 WR => WR2_IE,
		 CSR_WB_O => CSR_WB_O,
		 WB_O => WB_O,
		 BRANCH_O => SYNTHESIZED_WIRE_71,
		 ZERO_O => SYNTHESIZED_WIRE_106,
		 LESS_THAN_SIGNED_O => SYNTHESIZED_WIRE_107,
		 LESS_THAN_UNSIGNED_O => SYNTHESIZED_WIRE_108,
		 MEM_WR_O => MEM_WR_O,
		 FUNCT3_O => FUNCT3,
		 WR_O => WR_O);


b2v_inst59 : pip_reg_mem_wb
PORT MAP(CSR_WB => CSR_WB_O,
		 WB => WB_O,
		 CLK => CLK,
		 CLR => CLEAR,
		 WR => WR_O,
		 CSR_WB_O => SYNTHESIZED_WIRE_104,
		 WB_O => SYNTHESIZED_WIRE_109,
		 WR_O => SYNTHESIZED_WIRE_70);


b2v_inst6 : flag_reg
PORT MAP(FLAG_IN => EXP_INT_EN,
		 CLK => CLK,
		 CLR => CLEAR,
		 FLAG_OUT => EXP_INT_RETURN);


SYNTHESIZED_WIRE_53 <= WR_O(0) AND SYNTHESIZED_WIRE_95 AND SYNTHESIZED_WIRE_96;


SYNTHESIZED_WIRE_95 <= NOT(WR_O(1));



SYNTHESIZED_WIRE_96 <= NOT(WR_O(2));



b2v_inst8 : cla_32_add_1
PORT MAP(A => SYNTHESIZED_WIRE_100,
		 S => SYNTHESIZED_WIRE_101);


b2v_inst9 : alu
PORT MAP(DATAIN_1 => SYNTHESIZED_WIRE_98,
		 DATAIN_2 => SYNTHESIZED_WIRE_99,
		 OP => ALU_OP,
		 ZERO => SYNTHESIZED_WIRE_91,
		 LESS_THAN_SIGNED => SYNTHESIZED_WIRE_92,
		 LESS_THAN_UNSIGNED => SYNTHESIZED_WIRE_93,
		 DATA_OUT => SYNTHESIZED_WIRE_57);

PIN2_OUT <= EXP_PINS(0);
INT_EXTERNAL <= PIN1_IN;
PIN3_OUT <= EXP_PINS(1);
PIN4_OUT <= EXP_PINS(2);
PIN5_OUT <= EXP_PINS(3);

END bdf_type;